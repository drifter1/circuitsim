V1 5 0 2
V2 3 2 0.2
V3 7 6 2
R1 1 5 1.5
R2 1 12 1
R3 5 2 50
R4 5 6 0.1
R5 2 6 1.5
R6 3 4 0.2
R7 7 0 1e3
R8 4 0 10
I1 4 7 1e-3
I2 0 6 1e-3
C1 7 0 0.1
C2 2 0 0.2
L1 12 2 0.1
