R1 1 2 4
R2 2 0 2
V1 1 0 3
I1 0 2 2
